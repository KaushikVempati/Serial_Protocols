interface intf;
logic clk;
logic reset;
logic New_d;
logic rw_bar;
logic [6:0] Addr;
logic [7:0] Rdata;
logic [7:0] Wdata;
logic done_c;

logic SCLK_Ref;
 
endinterface
